NMOS Amplifier Circuit

*Model Declaration for NMOSFET
.model n NMOS W=10u L=0.5u VTO=1

*Gate Voltage for DC bias
Vgsq 1 0 dc 12

*Modulating Gate VOltage
Vgs 2 1 sin(0, 100m, 2000, 0, 0)
 
*Capacitor for decoupling
C1 2 3 50u

*Connection for NMOS
m1 4 3 0 0 n

*Drain Resistance
Rd 5 4 2.95k

*Voltage Divider
*Drain Gate
R1 5 3 329.15k
*Gate Source
R2 3 0 143.64k

*Drain Voltage
Vdd 5 0 dc 12

*Control Block
.control

*Transient Analysis Settings
tran 1us 2ms 

*File Write Setting
set appendwrite true
cd /Users/pushkalmishra/Desktop/Semester 3/Devices Lab/Experiment 9/NgSpice Code

*Command to write data
wrdata Amplifier_Circuit.txt v(2) - v(1)
wrdata Amplifier_Circuit.txt v(4)

.endc 