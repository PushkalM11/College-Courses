Half Wave Rectifier

*This code simulates a half wave bridge rectifier using
*A diode and a resistor

*Voltage Source-
V1 1 0 sin(0, 22, 50, 0, 0)

*Diode Model Declaration-
.model DMOD D

*Connection for Diode-
D1 1 2 DMOD

*Resistance connection-
R1 2 3 77.5

*Model for Battery
VDC 3 0 dc 12

*Control Block-
.control

*Transient Analysis Settings-
tran 1us 20ms

*Color Settings-
set color0 = white
set color1 = black
set color2 = blue

*Brushwidth Command-
set xbrushwidth = 3

*Plot Command for Voltage-
plot v(1) v(2) xlabel 'Time (in ms)' ylabel 'Voltage (in V)'

*Plot Command for Current-
plot i(VDC) xlabel 'Time (in ms)' ylabel 'Current (in mA)'

*Plot Command for Current and Voltage
plot v(2) 10*i(VDC) xlabel 'Time (in ms)'
    
.endc
