Full Wave Rectifier

*This code simulates a full wave bridge rectifier using
*Four diodes and a resistor

*Voltage Source-
V1 1 0 sin(0, 20, 50, 0, 0)

*Resistance connection-
R1 2 3 100

*Diode Components connection-
.model DMOD D

*Connection for Forward Bias-
D1 1 2 DMOD
D2 3 0 DMOD

*Connection for Reverse Bias-
D3 0 2 DMOD
D4 3 1 DMOD

*Model for Battery
VDC 2 3 dc 12

*Control Block-
.control

*Transient Analysis Settings-
tran 1ms 1s

*Color Settings-
set color0 = white
set color1 = black
set color2 = blue

*Plot Command for Voltage-
plot v(1) v(2)-V(3) xlabel 'Time (in s)' ylabel 'Voltage (in V)'

*Plot Command for Current-
plot i(VDC) xlabel 'Time (in s)' ylabel 'Current (in A)'
    
.endc
